library verilog;
use verilog.vl_types.all;
entity multiplier_tb is
end multiplier_tb;
