library verilog;
use verilog.vl_types.all;
entity MonPro_tb is
end MonPro_tb;
