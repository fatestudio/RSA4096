library verilog;
use verilog.vl_types.all;
entity file_readmemh_tb is
end file_readmemh_tb;
