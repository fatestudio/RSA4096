library verilog;
use verilog.vl_types.all;
entity ModExp_tb is
end ModExp_tb;
