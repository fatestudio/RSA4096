library verilog;
use verilog.vl_types.all;
entity MonExp_tb is
end MonExp_tb;
